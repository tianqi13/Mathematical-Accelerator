module mandelbrot_toplevel.sv(
    input logic rst,
    input logic clk,
    input logic en,
    input logic x_size,
    input logic y_size,
);

mapper MAPPER (

)

endmodule
