module ram_top(
    input logic clr,
    input logic enable,
    input logic clk,
    output logic 
);



endmodule
