module mandelbrot_toplevel.sv(

)

endmodule
